hello world how are things today
sample content
module dut
endmodule : dut
