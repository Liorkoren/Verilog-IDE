//module
module lior (ss, aa);
    output wire ss;
    input wire[31:0] aa;
endmodule