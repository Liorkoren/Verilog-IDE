module test #(parameter NO_DEFAULT) ();

endmodule