module generate_example();


  reg read,write = 0;

assign data_out = (read_v95) ? memory[address] : 0;

unrecognized statement;

reg [7:0] address1, address2;

assign data_out = (read_v95) ? memory[address] : 0;

endmodule;